module accumulator(rst, clk, out);

input rst, clk;
output [3:0] out;

// TODO

endmodule