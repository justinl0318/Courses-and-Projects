module baby_alu(in0, in1, alu_op, out);

input signed [7:0] in0, in1;
input [1:0] alu_op;
output reg signed [7:0] out;

// TODO

endmodule
